module not_gate(
    input logic a,
    output logic y
);

    
    assign y = ~a;

endmodule

